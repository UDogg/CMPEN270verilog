//Code an XOR gate using an "assign" statement
module xor_gate (output xor_Y, input xor_A, xor_B);
  assign xor_Y = xor_A ^ xor_B;   //complete this line
endmodule
