//Code an AND gate with an "assign" statement
module and_gate (output and_Y, input and_A, and_B);
  assign and_Y =and_A & and_B ;   //complete this line
endmodule
